module networking


struct Packet {
	packet_type u8
	data []u8
}


// Unsigned byte (0 to 255)
fn (mut p Packet) append_byte(value u8) {
	p.data = p.data.clone()
	p.data << value
}

// Signed byte (-128 to 127)
fn (mut p Packet) append_signed_byte(value i8) {
	p.data << u8(value)
}

// Signed fixed-point, 5 fractional bits (-4 to 3.96875)
fn (mut p Packet) append_signed_fixed_byte(value f32) {
	if value < -4.0 || value > 3.96875 {
		panic('Value out of range for signed fixed-point: $value')
	}

	p.data << u8((value + 4.0) * 32.0)
}

// Signed integer (-32768 to 32767)
fn (mut p Packet) append_short(value i16) {
	p.data << u8(value >> 8)
	p.data << u8(value & 0xFF)
}

// Signed fixed-point, 5 fractional bits (-1024 to 1023.96875)
fn (mut p Packet) append_signed_fixed_short(value f32) {
	if value < -1024.0 || value > 1023.96875 {
		panic('Value out of range for signed fixed-point: $value')
	}

	p.data << u8((value + 1024.0) * 32.0 >> 8)
	p.data << u8((value + 1024.0) * 32.0 & 0xFF)
}

// UTF-8 encoded string padded with spaces (0x20), length is always 64
fn (mut p Packet) append_string(value string) {
	if value.len > 64 {
		panic('String too long for packet: $value')
	}

	mut padded := value.bytes()
	padded << u8(0x20)

	for _ in padded.len .. 64 {
		padded << u8(0x20)
	}

	p.data << padded
}

// Binary data padded with null bytes (0x00) only if length is less than 1024
fn (mut p Packet) append_binary_data(value []u8) {
	if value.len > 1024 {
		panic('Binary data too long for packet: ${value.len} bytes')
	}

	mut padded := value.clone()
	for _ in padded.len .. 1024 {
		padded << u8(0x00)
	}

	p.data << padded
}


fn (mut p Packet) to_bytes() []u8 {
	mut bytes := []u8{len: 1 + p.data.len}
	bytes[0] = p.packet_type

	if p.data.len > 0 {
		bytes[1..] = p.data
	}

	return bytes
}